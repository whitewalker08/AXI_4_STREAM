class ei_AXIS_coverage_packet;
  int sparse_stream;
  int aligned_stream;
  int unaligned_stream;
  int num_trans;
  bit TLAST;  
endclass : ei_AXIS_coverage_packet
