/*-----------------------------------------------------------------------------



File name    : ei_AXIS_include_all.svh



Title        : AXI_stream_include_all_file



Project      : AXIS_SV_VIP  



Created On   : 02-06-2022



Developers   : einfochips Ltd



Purpose      : to include all file in one single file and use them in testbench file.

               
-------------------------------------------------------------------------------

Copyright (c) 2000-2006 eInfochips           - All rights reserved



This software is authored by eInfochips and is eInfochips intellectual

property, including the copyrights in all countries in the world. This

software is provided under a license to use only with all other rights,

including ownership rights, being retained by eInfochips



This file may not be distributed, copied, or reproduced in any manner,

electronic or otherwise, without the express written consent of

eInfochips

-------------------------------------------------------------------------------

Revision: 1.0

-------------------------------------------------------------------------------*/
`include "ei_AXIS_config.sv"
`include "ei_AXIS_master_interface.sv"
`include "ei_AXIS_slave_interface.sv"
`include "ei_AXIS_interconnect.sv"
`include "ei_AXIS_master_transaction.sv"
`include "ei_AXIS_master_generator.sv"
`include "ei_AXIS_master_driver.sv"
`include "ei_AXIS_coverage_packet.sv"
`include "ei_AXIS_master_monitor.sv"
`include "ei_AXIS_coverage.sv"
`include "ei_AXIS_slave_driver.sv"
`include "ei_AXIS_slave_monitor.sv"
`include "ei_AXIS_scoreboard.sv"
`include "ei_AXIS_master_agent.sv"
`include "ei_AXIS_slave_agent.sv"
`include "ei_AXIS_environment.sv"
`include "ei_AXIS_write.sv"
`include "ei_AXIS_unaligned_stream.sv"
`include "ei_AXIS_sparse_stream.sv"
`include "ei_AXIS_single_transfer_with_pos.sv"
`include "ei_AXIS_aligned_sparse.sv"
`include "ei_AXIS_aligned_unaligned.sv"
`include "ei_AXIS_sparse_unaligned.sv"
`include "ei_AXIS_sparse_aligned_unaligned.sv"
`include "ei_AXIS_video_frame.sv"
`include "ei_AXIS_test.sv"


/*-------------------------------------------------------------------------------

Copyright (c) 2000-2006 eInfochips           - All rights reserved



This software is authored by eInfochips and is eInfochips intellectual

property, including the copyrights in all countries in the world. This

software is provided under a license to use only with all other rights,

including ownership rights, being retained by eInfochips



This file may not be distributed, copied, or reproduced in any manner,

electronic or otherwise, without the express written consent of

eInfochips

-------------------------------------------------------------------------------

Revision: 1.0

-------------------------------------------------------------------------------*/
